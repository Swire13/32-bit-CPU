`timescale 1ns/1ps

module CPU_TB ();

reg CLK_DUT = 1'b0;
reg RST_DUT;
reg [31:0] DATA_IN_DUT;
reg [31:0] INSTR_IN_DUT;
wire [31:0] DATA_OUT_DUT;
wire [31:0] DADDR_DUT;
wire DWR_DUT;
wire DEN_DUT;
wire [31:0] IADDR_DUT;
wire IEN_DUT;

reg [31:0] data[0:255];
reg [31:0] instr[0:255];
integer i;

CPU DUT(
  .clk (CLK_DUT),
  .RST (RST_DUT),
  .DATA_IN (DATA_IN_DUT),
  .INSTR_IN (INSTR_IN_DUT),
  .DATA_OUT (DATA_OUT_DUT),
  .DADDR (DADDR_DUT),
  .DWR (DWR_DUT),
  .DEN (DEN_DUT),
  .IADDR (IADDR_DUT),
  .IEN (IEN_DUT)
);

initial begin
   for (i = 0; i < 256; i = i + 1) begin
     data[i] = 32'b00000000000000000000000000000000;
   end
   instr[0]  = 32'b1_0000000000000000000000000000011;//JMP
   instr[1]  = 32'b00000000000000000000000000000000;//NOP
   instr[2]  = 32'b00000000000000000000000000000000;//NOP
   instr[3]  = 32'b01_000000000000_000000_000001100100;//LD    R0 = 100
   instr[4]  = 32'b01_000000000000_000001_000000001010;//LD    R1 = 10
   instr[5]  = 32'b01_000000000000_111111_000000000110;//LD    R63 = 6
   instr[6]  = 32'b0000010_0000000_000000_000001_000000;//SUB  R0 = R0 - R1
   instr[7]  = 32'b0011_0000000000000000_111111_000000;//BNE
   instr[8]  = 32'b01_000000000010_000101_010001101101;//LD    R5 = 1133
   instr[9]  = 32'b01_000000000000_111110_000000000000;//LD    R62 = 0
   instr[10]  = 32'b00010_000000000000000_111110_000101;//WR   MEM[R62] = R5
   instr[11]  = 32'b00011_000000000_000110_111110_000000;//RD  R6 = MEM[R62]
   instr[12]  = 32'b01_000000000000_111101_000000001111;//LD   R61 = 15
   instr[13]  = 32'b0010_0010010001101101_111101_000110;//BEQ  
   instr[14]  = 32'b00000000000000000000000000000000;//NOP
   instr[15]  = 32'b00000000000000000000000000000000;//NOP
   instr[16]  = 32'b01_111010100000_000000_010011011010;//LD    R0 = 15336666
   instr[17]  = 32'b01_000000000000_000001_000010011011;//LD    R1 = 155
   instr[18]  = 32'b0000001_0000000_000010_000001_000000;//ADD  R2 = R0 + R1
   instr[19]  = 32'b0000010_0000000_000011_000001_000000;//SUB  R3 = R0 - R1
   instr[20]  = 32'b0000011_0000000_000100_000001_000000;//AND  R4 = R0 & R1
   instr[21]  = 32'b0000100_0000000_000101_000001_000000;//OR   R5 = R0 | R1
   instr[22]  = 32'b0000101_0000000_000110_000001_000000;//XOR  R6 = R0 ^ R1
   instr[23]  = 32'b0000110_0000000_000111_000001_0_00101;//SHL R7 = R0 << 5
   instr[24]  = 32'b0000110_0000000_001000_000001_1_11010;//ROL R8 = R1 <<< 26
   instr[25]  = 32'b0000111_0000000_001001_000001_0_00100;//SHR R9 = R0 >> 4
   instr[26]  = 32'b0000111_0000000_001010_000001_1_00011;//ROR R10 = R1 >>> 3
   instr[27]  = 32'b01_000000000000_001011_000000000000;//LD    
   instr[28]  = 32'b01_000000000000_001100_000000000001;//LD
   instr[29]  = 32'b01_000000000000_001101_000000000010;//LD
   instr[30]  = 32'b01_000000000000_001110_000000000011;//LD
   instr[31]  = 32'b01_000000000000_001111_000000000100;//LD
   instr[32]  = 32'b01_000000000000_010000_000000000101;//LD
   instr[33]  = 32'b01_000000000000_010001_000000000110;//LD
   instr[34]  = 32'b01_000000000000_010010_000000000111;//LD
   instr[35]  = 32'b01_000000000000_010011_000000001000;//LD
   instr[36]  = 32'b01_000000000000_010100_000000001001;//LD
   instr[37]  = 32'b01_000000000000_010101_000000001010;//LD
   instr[38]  = 32'b00010_000000000000000_001011_000010;//WR
   instr[39]  = 32'b00010_000000000000000_001100_000011;//WR
   instr[40]  = 32'b00010_000000000000000_001101_000100;//WR
   instr[41]  = 32'b00010_000000000000000_001110_000101;//WR
   instr[42]  = 32'b00010_000000000000000_001111_000110;//WR
   instr[43]  = 32'b00010_000000000000000_010000_000111;//WR
   instr[44]  = 32'b00010_000000000000000_010001_001000;//WR
   instr[45]  = 32'b00010_000000000000000_010010_001001;//WR
   instr[46]  = 32'b00010_000000000000000_010011_001010;//WR
   instr[47]  = 32'b00010_000000000000000_010100_001011;//WR
   instr[48]  = 32'b00010_000000000000000_010101_001100;//WR
   for (i = 49; i < 256; i = i + 1) begin
     data[i] = 32'b1_0000000000000000000000000000000;//JMP
   end
   RST_DUT = 1'b1;
	#12;
	RST_DUT = 1'b0;
	#480;
	for (i = 0; i < 256; i = i + 1) 
     $display("data[%d]: %b", i, data[i]);
end

always @(posedge CLK_DUT) begin
  INSTR_IN_DUT <= instr[IADDR_DUT];
end	

always @(posedge CLK_DUT) begin
  if (DEN_DUT == 1'b1) begin
	 if (DWR_DUT == 1'b1)
		data[DADDR_DUT] = DATA_OUT_DUT;
	 else
		DATA_IN_DUT = data[DADDR_DUT];
  end	else begin
    DATA_IN_DUT <= 32'h00000000;
  end
end

always #5 CLK_DUT = ~CLK_DUT;

endmodule